//header guards
`ifndef _registerFile_vh_
`define _registerFile_vh_

`include "decoders.v"
`include "tristate.v"
`include "DFFwithEnable.v"

/*Note: The register FILE outputs/changes RD DATAs as soon as RD ADDRESSes are changed
Doesn't wait for clock | may need to introduce DFF for read ADDRESSES*/

module registers(RDADDRESS1,RDADDRESS2,WRADDRESS,WRDATA,read,write,RDOUT1,RDOUT2,clk);

	input[4:0] RDADDRESS1,RDADDRESS2,WRADDRESS;
	input[31:0] WRDATA;

	input read,write,clk;

	output[31:0] RDOUT1,RDOUT2;

	//module decoder5x32(enable,IN,OUT);
	wire[31:0] WRDECODER_OUT;
	decoder5x32 WRDecoder(write,WRADDRESS,WRDECODER_OUT);

	wire[31:0] DFF_OUT[0:31];
	//module DFF32bitEnable(DATAIN,clk,DATAOUT,load);

	//WRITE DATA into REGISTER FILE
	DFF32bitEnable DFF0(WRDATA,clk,DFF_OUT[0],WRDECODER_OUT[0]);
	DFF32bitEnable DFF1(WRDATA,clk,DFF_OUT[1],WRDECODER_OUT[1]);
	DFF32bitEnable DFF2(WRDATA,clk,DFF_OUT[2],WRDECODER_OUT[2]);
	DFF32bitEnable DFF3(WRDATA,clk,DFF_OUT[3],WRDECODER_OUT[3]);
	DFF32bitEnable DFF4(WRDATA,clk,DFF_OUT[4],WRDECODER_OUT[4]);
	DFF32bitEnable DFF5(WRDATA,clk,DFF_OUT[5],WRDECODER_OUT[5]);
	DFF32bitEnable DFF6(WRDATA,clk,DFF_OUT[6],WRDECODER_OUT[6]);
	DFF32bitEnable DFF7(WRDATA,clk,DFF_OUT[7],WRDECODER_OUT[7]);
	DFF32bitEnable DFF8(WRDATA,clk,DFF_OUT[8],WRDECODER_OUT[8]);
	DFF32bitEnable DFF9(WRDATA,clk,DFF_OUT[9],WRDECODER_OUT[9]);
	DFF32bitEnable DFF10(WRDATA,clk,DFF_OUT[10],WRDECODER_OUT[10]);
	DFF32bitEnable DFF11(WRDATA,clk,DFF_OUT[11],WRDECODER_OUT[11]);
	DFF32bitEnable DFF12(WRDATA,clk,DFF_OUT[12],WRDECODER_OUT[12]);
	DFF32bitEnable DFF13(WRDATA,clk,DFF_OUT[13],WRDECODER_OUT[13]);
	DFF32bitEnable DFF14(WRDATA,clk,DFF_OUT[14],WRDECODER_OUT[14]);
	DFF32bitEnable DFF15(WRDATA,clk,DFF_OUT[15],WRDECODER_OUT[15]);
	DFF32bitEnable DFF16(WRDATA,clk,DFF_OUT[16],WRDECODER_OUT[16]);
	DFF32bitEnable DFF17(WRDATA,clk,DFF_OUT[17],WRDECODER_OUT[17]);
	DFF32bitEnable DFF18(WRDATA,clk,DFF_OUT[18],WRDECODER_OUT[18]);
	DFF32bitEnable DFF19(WRDATA,clk,DFF_OUT[19],WRDECODER_OUT[19]);
	DFF32bitEnable DFF20(WRDATA,clk,DFF_OUT[20],WRDECODER_OUT[20]);
	DFF32bitEnable DFF21(WRDATA,clk,DFF_OUT[21],WRDECODER_OUT[21]);
	DFF32bitEnable DFF22(WRDATA,clk,DFF_OUT[22],WRDECODER_OUT[22]);
	DFF32bitEnable DFF23(WRDATA,clk,DFF_OUT[23],WRDECODER_OUT[23]);
	DFF32bitEnable DFF24(WRDATA,clk,DFF_OUT[24],WRDECODER_OUT[24]);
	DFF32bitEnable DFF25(WRDATA,clk,DFF_OUT[25],WRDECODER_OUT[25]);
	DFF32bitEnable DFF26(WRDATA,clk,DFF_OUT[26],WRDECODER_OUT[26]);
	DFF32bitEnable DFF27(WRDATA,clk,DFF_OUT[27],WRDECODER_OUT[27]);
	DFF32bitEnable DFF28(WRDATA,clk,DFF_OUT[28],WRDECODER_OUT[28]);
	DFF32bitEnable DFF29(WRDATA,clk,DFF_OUT[29],WRDECODER_OUT[29]);
	DFF32bitEnable DFF30(WRDATA,clk,DFF_OUT[30],WRDECODER_OUT[30]);
	DFF32bitEnable DFF31(WRDATA,clk,DFF_OUT[31],WRDECODER_OUT[31]);


	//READ DATA from REGISTER FILE
	wire[31:0] RD1DECODER_OUT,RD2DECODER_OUT;

	//module decoder5x32(enable,IN,OUT);
	decoder5x32 RD1Decoder(read,RDADDRESS1,RD1DECODER_OUT);
	decoder5x32 RD2Decoder(read,RDADDRESS2,RD2DECODER_OUT);

	//module tristate32bit (DATAIN,enable,DATAOUT);
	tristate32bit DFF0_RD1OUT(DFF_OUT[0],RD1DECODER_OUT[0],RDOUT1);
	tristate32bit DFF1_RD1OUT(DFF_OUT[1],RD1DECODER_OUT[1],RDOUT1);
	tristate32bit DFF2_RD1OUT(DFF_OUT[2],RD1DECODER_OUT[2],RDOUT1);
	tristate32bit DFF3_RD1OUT(DFF_OUT[3],RD1DECODER_OUT[3],RDOUT1);
	tristate32bit DFF4_RD1OUT(DFF_OUT[4],RD1DECODER_OUT[4],RDOUT1);
	tristate32bit DFF5_RD1OUT(DFF_OUT[5],RD1DECODER_OUT[5],RDOUT1);
	tristate32bit DFF6_RD1OUT(DFF_OUT[6],RD1DECODER_OUT[6],RDOUT1);
	tristate32bit DFF7_RD1OUT(DFF_OUT[7],RD1DECODER_OUT[7],RDOUT1);
	tristate32bit DFF8_RD1OUT(DFF_OUT[8],RD1DECODER_OUT[8],RDOUT1);
	tristate32bit DFF9_RD1OUT(DFF_OUT[9],RD1DECODER_OUT[9],RDOUT1);
	tristate32bit DFF10_RD1OUT(DFF_OUT[10],RD1DECODER_OUT[10],RDOUT1);
	tristate32bit DFF11_RD1OUT(DFF_OUT[11],RD1DECODER_OUT[11],RDOUT1);
	tristate32bit DFF12_RD1OUT(DFF_OUT[12],RD1DECODER_OUT[12],RDOUT1);
	tristate32bit DFF13_RD1OUT(DFF_OUT[13],RD1DECODER_OUT[13],RDOUT1);
	tristate32bit DFF14_RD1OUT(DFF_OUT[14],RD1DECODER_OUT[14],RDOUT1);
	tristate32bit DFF15_RD1OUT(DFF_OUT[15],RD1DECODER_OUT[15],RDOUT1);
	tristate32bit DFF16_RD1OUT(DFF_OUT[16],RD1DECODER_OUT[16],RDOUT1);
	tristate32bit DFF17_RD1OUT(DFF_OUT[17],RD1DECODER_OUT[17],RDOUT1);
	tristate32bit DFF18_RD1OUT(DFF_OUT[18],RD1DECODER_OUT[18],RDOUT1);
	tristate32bit DFF19_RD1OUT(DFF_OUT[19],RD1DECODER_OUT[19],RDOUT1);
	tristate32bit DFF20_RD1OUT(DFF_OUT[20],RD1DECODER_OUT[20],RDOUT1);
	tristate32bit DFF21_RD1OUT(DFF_OUT[21],RD1DECODER_OUT[21],RDOUT1);
	tristate32bit DFF22_RD1OUT(DFF_OUT[22],RD1DECODER_OUT[22],RDOUT1);
	tristate32bit DFF23_RD1OUT(DFF_OUT[23],RD1DECODER_OUT[23],RDOUT1);
	tristate32bit DFF24_RD1OUT(DFF_OUT[24],RD1DECODER_OUT[24],RDOUT1);
	tristate32bit DFF25_RD1OUT(DFF_OUT[25],RD1DECODER_OUT[25],RDOUT1);
	tristate32bit DFF26_RD1OUT(DFF_OUT[26],RD1DECODER_OUT[26],RDOUT1);
	tristate32bit DFF27_RD1OUT(DFF_OUT[27],RD1DECODER_OUT[27],RDOUT1);
	tristate32bit DFF28_RD1OUT(DFF_OUT[28],RD1DECODER_OUT[28],RDOUT1);
	tristate32bit DFF29_RD1OUT(DFF_OUT[29],RD1DECODER_OUT[29],RDOUT1);
	tristate32bit DFF30_RD1OUT(DFF_OUT[30],RD1DECODER_OUT[30],RDOUT1);
	tristate32bit DFF31_RD1OUT(DFF_OUT[31],RD1DECODER_OUT[31],RDOUT1);


	tristate32bit DFF0_RD2OUT(DFF_OUT[0],RD2DECODER_OUT[0],RDOUT2);
	tristate32bit DFF1_RD2OUT(DFF_OUT[1],RD2DECODER_OUT[1],RDOUT2);
	tristate32bit DFF2_RD2OUT(DFF_OUT[2],RD2DECODER_OUT[2],RDOUT2);
	tristate32bit DFF3_RD2OUT(DFF_OUT[3],RD2DECODER_OUT[3],RDOUT2);
	tristate32bit DFF4_RD2OUT(DFF_OUT[4],RD2DECODER_OUT[4],RDOUT2);
	tristate32bit DFF5_RD2OUT(DFF_OUT[5],RD2DECODER_OUT[5],RDOUT2);
	tristate32bit DFF6_RD2OUT(DFF_OUT[6],RD2DECODER_OUT[6],RDOUT2);
	tristate32bit DFF7_RD2OUT(DFF_OUT[7],RD2DECODER_OUT[7],RDOUT2);
	tristate32bit DFF8_RD2OUT(DFF_OUT[8],RD2DECODER_OUT[8],RDOUT2);
	tristate32bit DFF9_RD2OUT(DFF_OUT[9],RD2DECODER_OUT[9],RDOUT2);
	tristate32bit DFF10_RD2OUT(DFF_OUT[10],RD2DECODER_OUT[10],RDOUT2);
	tristate32bit DFF11_RD2OUT(DFF_OUT[11],RD2DECODER_OUT[11],RDOUT2);
	tristate32bit DFF12_RD2OUT(DFF_OUT[12],RD2DECODER_OUT[12],RDOUT2);
	tristate32bit DFF13_RD2OUT(DFF_OUT[13],RD2DECODER_OUT[13],RDOUT2);
	tristate32bit DFF14_RD2OUT(DFF_OUT[14],RD2DECODER_OUT[14],RDOUT2);
	tristate32bit DFF15_RD2OUT(DFF_OUT[15],RD2DECODER_OUT[15],RDOUT2);
	tristate32bit DFF16_RD2OUT(DFF_OUT[16],RD2DECODER_OUT[16],RDOUT2);
	tristate32bit DFF17_RD2OUT(DFF_OUT[17],RD2DECODER_OUT[17],RDOUT2);
	tristate32bit DFF18_RD2OUT(DFF_OUT[18],RD2DECODER_OUT[18],RDOUT2);
	tristate32bit DFF19_RD2OUT(DFF_OUT[19],RD2DECODER_OUT[19],RDOUT2);
	tristate32bit DFF20_RD2OUT(DFF_OUT[20],RD2DECODER_OUT[20],RDOUT2);
	tristate32bit DFF21_RD2OUT(DFF_OUT[21],RD2DECODER_OUT[21],RDOUT2);
	tristate32bit DFF22_RD2OUT(DFF_OUT[22],RD2DECODER_OUT[22],RDOUT2);
	tristate32bit DFF23_RD2OUT(DFF_OUT[23],RD2DECODER_OUT[23],RDOUT2);
	tristate32bit DFF24_RD2OUT(DFF_OUT[24],RD2DECODER_OUT[24],RDOUT2);
	tristate32bit DFF25_RD2OUT(DFF_OUT[25],RD2DECODER_OUT[25],RDOUT2);
	tristate32bit DFF26_RD2OUT(DFF_OUT[26],RD2DECODER_OUT[26],RDOUT2);
	tristate32bit DFF27_RD2OUT(DFF_OUT[27],RD2DECODER_OUT[27],RDOUT2);
	tristate32bit DFF28_RD2OUT(DFF_OUT[28],RD2DECODER_OUT[28],RDOUT2);
	tristate32bit DFF29_RD2OUT(DFF_OUT[29],RD2DECODER_OUT[29],RDOUT2);
	tristate32bit DFF30_RD2OUT(DFF_OUT[30],RD2DECODER_OUT[30],RDOUT2);
	tristate32bit DFF31_RD2OUT(DFF_OUT[31],RD2DECODER_OUT[31],RDOUT2);

endmodule // registers

`endif
