//header guards
`ifndef _MUX_all_vh_
`define _MUX_all_vh_

`include "D-FlipFlop.v"

module MUX_2x1(A,select,out);
	input[1:0] A;
	input select;

	output out;

	assign out=A[0]&(~select)|A[1]&select;

endmodule

//2x1 MUX 
module MUX2x1(data0,data1,select,out);
	input data0,data1,select;
	output out;
	
	assign out = data0 & (~select) | data1 & select;

endmodule // MUX2x1

module MUX8bit_2x1(DATA0,DATA1,select,OUT);

	input[7:0] DATA0, DATA1;
	input select;

	output[7:0] OUT;

	MUX2x1 MUX0(DATA0[0],DATA1[0],select,OUT[0]);
	MUX2x1 MUX1(DATA0[1],DATA1[1],select,OUT[1]);
	MUX2x1 MUX2(DATA0[2],DATA1[2],select,OUT[2]);
	MUX2x1 MUX3(DATA0[3],DATA1[3],select,OUT[3]);
	MUX2x1 MUX4(DATA0[4],DATA1[4],select,OUT[4]);
	MUX2x1 MUX5(DATA0[5],DATA1[5],select,OUT[5]);
	MUX2x1 MUX6(DATA0[6],DATA1[6],select,OUT[6]);
	MUX2x1 MUX7(DATA0[7],DATA1[7],select,OUT[7]);

endmodule //MUX8bit_2x1


module MUX24bit_2x1(DATA0,DATA1,select,OUT);

	input[23:0] DATA0,DATA1;
	input select;

	output[23:0] OUT;

  //MUX2x1 MUX0(DATA0[0],DATA1[0],select,OUT[0]);
	MUX2x1 MUX0(DATA0[0],DATA1[0],select,OUT[0]);
	MUX2x1 MUX1(DATA0[1],DATA1[1],select,OUT[1]);
	MUX2x1 MUX2(DATA0[2],DATA1[2],select,OUT[2]);
	MUX2x1 MUX3(DATA0[3],DATA1[3],select,OUT[3]);
	MUX2x1 MUX4(DATA0[4],DATA1[4],select,OUT[4]);
	MUX2x1 MUX5(DATA0[5],DATA1[5],select,OUT[5]);
	MUX2x1 MUX6(DATA0[6],DATA1[6],select,OUT[6]);
	MUX2x1 MUX7(DATA0[7],DATA1[7],select,OUT[7]);
	MUX2x1 MUX8(DATA0[8],DATA1[8],select,OUT[8]);
	MUX2x1 MUX9(DATA0[9],DATA1[9],select,OUT[9]);
	MUX2x1 MUX10(DATA0[10],DATA1[10],select,OUT[10]);
	MUX2x1 MUX11(DATA0[11],DATA1[11],select,OUT[11]);
	MUX2x1 MUX12(DATA0[12],DATA1[12],select,OUT[12]);
	MUX2x1 MUX13(DATA0[13],DATA1[13],select,OUT[13]);
	MUX2x1 MUX14(DATA0[14],DATA1[14],select,OUT[14]);
	MUX2x1 MUX15(DATA0[15],DATA1[15],select,OUT[15]);
	MUX2x1 MUX16(DATA0[16],DATA1[16],select,OUT[16]);
	MUX2x1 MUX17(DATA0[17],DATA1[17],select,OUT[17]);
	MUX2x1 MUX18(DATA0[18],DATA1[18],select,OUT[18]);
	MUX2x1 MUX19(DATA0[19],DATA1[19],select,OUT[19]);
	MUX2x1 MUX20(DATA0[20],DATA1[20],select,OUT[20]);
	MUX2x1 MUX21(DATA0[21],DATA1[21],select,OUT[21]);
	MUX2x1 MUX22(DATA0[22],DATA1[22],select,OUT[22]);
	MUX2x1 MUX23(DATA0[23],DATA1[23],select,OUT[23]);
	
endmodule // MUX24bit_2x1


module MUX32bit_2x1(DATA0,DATA1,select,OUT);

	input[31:0] DATA0,DATA1;
	input select;

	output[31:0] OUT;

  //MUX2x1 MUX0(DATA0[0],DATA1[0],select,OUT[0]);
	MUX2x1 MUX0(DATA0[0],DATA1[0],select,OUT[0]);
	MUX2x1 MUX1(DATA0[1],DATA1[1],select,OUT[1]);
	MUX2x1 MUX2(DATA0[2],DATA1[2],select,OUT[2]);
	MUX2x1 MUX3(DATA0[3],DATA1[3],select,OUT[3]);
	MUX2x1 MUX4(DATA0[4],DATA1[4],select,OUT[4]);
	MUX2x1 MUX5(DATA0[5],DATA1[5],select,OUT[5]);
	MUX2x1 MUX6(DATA0[6],DATA1[6],select,OUT[6]);
	MUX2x1 MUX7(DATA0[7],DATA1[7],select,OUT[7]);
	MUX2x1 MUX8(DATA0[8],DATA1[8],select,OUT[8]);
	MUX2x1 MUX9(DATA0[9],DATA1[9],select,OUT[9]);
	MUX2x1 MUX10(DATA0[10],DATA1[10],select,OUT[10]);
	MUX2x1 MUX11(DATA0[11],DATA1[11],select,OUT[11]);
	MUX2x1 MUX12(DATA0[12],DATA1[12],select,OUT[12]);
	MUX2x1 MUX13(DATA0[13],DATA1[13],select,OUT[13]);
	MUX2x1 MUX14(DATA0[14],DATA1[14],select,OUT[14]);
	MUX2x1 MUX15(DATA0[15],DATA1[15],select,OUT[15]);
	MUX2x1 MUX16(DATA0[16],DATA1[16],select,OUT[16]);
	MUX2x1 MUX17(DATA0[17],DATA1[17],select,OUT[17]);
	MUX2x1 MUX18(DATA0[18],DATA1[18],select,OUT[18]);
	MUX2x1 MUX19(DATA0[19],DATA1[19],select,OUT[19]);
	MUX2x1 MUX20(DATA0[20],DATA1[20],select,OUT[20]);
	MUX2x1 MUX21(DATA0[21],DATA1[21],select,OUT[21]);
	MUX2x1 MUX22(DATA0[22],DATA1[22],select,OUT[22]);
	MUX2x1 MUX23(DATA0[23],DATA1[23],select,OUT[23]);
	MUX2x1 MUX24(DATA0[24],DATA1[24],select,OUT[24]);
	MUX2x1 MUX25(DATA0[25],DATA1[25],select,OUT[25]);
	MUX2x1 MUX26(DATA0[26],DATA1[26],select,OUT[26]);
	MUX2x1 MUX27(DATA0[27],DATA1[27],select,OUT[27]);
	MUX2x1 MUX28(DATA0[28],DATA1[28],select,OUT[28]);
	MUX2x1 MUX29(DATA0[29],DATA1[29],select,OUT[29]);
	MUX2x1 MUX30(DATA0[30],DATA1[30],select,OUT[30]);
	MUX2x1 MUX31(DATA0[31],DATA1[31],select,OUT[31]);
endmodule // MUX32bit_2x1


//Right shift by 1 unit, if shift=1
//for use in FPM
module MUX_24bitShifter(DATA,shift,OUT);

	input[23:0] DATA;
	input shift;

	output[23:0] OUT;

	MUX2x1 MUX0(DATA[0],DATA[1],shift,OUT[0]);
	MUX2x1 MUX1(DATA[1],DATA[2],shift,OUT[1]);
	MUX2x1 MUX2(DATA[2],DATA[3],shift,OUT[2]);
	MUX2x1 MUX3(DATA[3],DATA[4],shift,OUT[3]);
	MUX2x1 MUX4(DATA[4],DATA[5],shift,OUT[4]);
	MUX2x1 MUX5(DATA[5],DATA[6],shift,OUT[5]);
	MUX2x1 MUX6(DATA[6],DATA[7],shift,OUT[6]);
	MUX2x1 MUX7(DATA[7],DATA[8],shift,OUT[7]);
	MUX2x1 MUX8(DATA[8],DATA[9],shift,OUT[8]);
	MUX2x1 MUX9(DATA[9],DATA[10],shift,OUT[9]);
	MUX2x1 MUX10(DATA[10],DATA[11],shift,OUT[10]);
	MUX2x1 MUX11(DATA[11],DATA[12],shift,OUT[11]);
	MUX2x1 MUX12(DATA[12],DATA[13],shift,OUT[12]);
	MUX2x1 MUX13(DATA[13],DATA[14],shift,OUT[13]);
	MUX2x1 MUX14(DATA[14],DATA[15],shift,OUT[14]);
	MUX2x1 MUX15(DATA[15],DATA[16],shift,OUT[15]);
	MUX2x1 MUX16(DATA[16],DATA[17],shift,OUT[16]);
	MUX2x1 MUX17(DATA[17],DATA[18],shift,OUT[17]);
	MUX2x1 MUX18(DATA[18],DATA[19],shift,OUT[18]);
	MUX2x1 MUX19(DATA[19],DATA[20],shift,OUT[19]);
	MUX2x1 MUX20(DATA[20],DATA[21],shift,OUT[20]);
	MUX2x1 MUX21(DATA[21],DATA[22],shift,OUT[21]);
	MUX2x1 MUX22(DATA[22],DATA[23],shift,OUT[22]);
	MUX2x1 MUX23(DATA[23],0,shift,OUT[23]);

endmodule

//2x1 MUX with D-Flip Flop(with clock) at OUTPUT
//for use in Barrel Shifter
module MUX2x1_DFF(data0,data1,select,out,clk);
	input data0,data1,select,clk;
	output out;

	wire mux_out;

	assign mux_out = data0 & (~select) | data1 & select;
	DFlipFlop DFF(mux_out,clk,out);

endmodule // MUX2x1_DFF


module MUX4x1(data0,data1,data2,data3,SELECT,out,clk);

	input data0,data1,data2,data3,clk;
	input[1:0] SELECT;

	output out;

	wire level1_MUX0_out,level1_MUX1_out;
	MUX2x1 level1_MUX0(data0,data1,SELECT[0],level1_MUX0_out);
	MUX2x1 level1_MUX1(data2,data3,SELECT[0],level1_MUX1_out);

	MUX2x1 level2_MUX(level1_MUX0_out,level1_MUX1_out,SELECT[1],out);
endmodule // MUX4x1


module MUX64bit_4x1(DATA0,DATA1,DATA2,DATA3,SELECT,OUT,clk);

	input[63:0] DATA0,DATA1,DATA2,DATA3;
	input[1:0] SELECT;
	input clk;

	output[63:0] OUT;

	MUX4x1 MUX0(DATA0[0],DATA1[0],DATA2[0],DATA3[0],SELECT,OUT[0],clk);
	MUX4x1 MUX1(DATA0[1],DATA1[1],DATA2[1],DATA3[1],SELECT,OUT[1],clk);
	MUX4x1 MUX2(DATA0[2],DATA1[2],DATA2[2],DATA3[2],SELECT,OUT[2],clk);
	MUX4x1 MUX3(DATA0[3],DATA1[3],DATA2[3],DATA3[3],SELECT,OUT[3],clk);
	MUX4x1 MUX4(DATA0[4],DATA1[4],DATA2[4],DATA3[4],SELECT,OUT[4],clk);
	MUX4x1 MUX5(DATA0[5],DATA1[5],DATA2[5],DATA3[5],SELECT,OUT[5],clk);
	MUX4x1 MUX6(DATA0[6],DATA1[6],DATA2[6],DATA3[6],SELECT,OUT[6],clk);
	MUX4x1 MUX7(DATA0[7],DATA1[7],DATA2[7],DATA3[7],SELECT,OUT[7],clk);
	MUX4x1 MUX8(DATA0[8],DATA1[8],DATA2[8],DATA3[8],SELECT,OUT[8],clk);
	MUX4x1 MUX9(DATA0[9],DATA1[9],DATA2[9],DATA3[9],SELECT,OUT[9],clk);
	MUX4x1 MUX10(DATA0[10],DATA1[10],DATA2[10],DATA3[10],SELECT,OUT[10],clk);
	MUX4x1 MUX11(DATA0[11],DATA1[11],DATA2[11],DATA3[11],SELECT,OUT[11],clk);
	MUX4x1 MUX12(DATA0[12],DATA1[12],DATA2[12],DATA3[12],SELECT,OUT[12],clk);
	MUX4x1 MUX13(DATA0[13],DATA1[13],DATA2[13],DATA3[13],SELECT,OUT[13],clk);
	MUX4x1 MUX14(DATA0[14],DATA1[14],DATA2[14],DATA3[14],SELECT,OUT[14],clk);
	MUX4x1 MUX15(DATA0[15],DATA1[15],DATA2[15],DATA3[15],SELECT,OUT[15],clk);
	MUX4x1 MUX16(DATA0[16],DATA1[16],DATA2[16],DATA3[16],SELECT,OUT[16],clk);
	MUX4x1 MUX17(DATA0[17],DATA1[17],DATA2[17],DATA3[17],SELECT,OUT[17],clk);
	MUX4x1 MUX18(DATA0[18],DATA1[18],DATA2[18],DATA3[18],SELECT,OUT[18],clk);
	MUX4x1 MUX19(DATA0[19],DATA1[19],DATA2[19],DATA3[19],SELECT,OUT[19],clk);
	MUX4x1 MUX20(DATA0[20],DATA1[20],DATA2[20],DATA3[20],SELECT,OUT[20],clk);
	MUX4x1 MUX21(DATA0[21],DATA1[21],DATA2[21],DATA3[21],SELECT,OUT[21],clk);
	MUX4x1 MUX22(DATA0[22],DATA1[22],DATA2[22],DATA3[22],SELECT,OUT[22],clk);
	MUX4x1 MUX23(DATA0[23],DATA1[23],DATA2[23],DATA3[23],SELECT,OUT[23],clk);
	MUX4x1 MUX24(DATA0[24],DATA1[24],DATA2[24],DATA3[24],SELECT,OUT[24],clk);
	MUX4x1 MUX25(DATA0[25],DATA1[25],DATA2[25],DATA3[25],SELECT,OUT[25],clk);
	MUX4x1 MUX26(DATA0[26],DATA1[26],DATA2[26],DATA3[26],SELECT,OUT[26],clk);
	MUX4x1 MUX27(DATA0[27],DATA1[27],DATA2[27],DATA3[27],SELECT,OUT[27],clk);
	MUX4x1 MUX28(DATA0[28],DATA1[28],DATA2[28],DATA3[28],SELECT,OUT[28],clk);
	MUX4x1 MUX29(DATA0[29],DATA1[29],DATA2[29],DATA3[29],SELECT,OUT[29],clk);
	MUX4x1 MUX30(DATA0[30],DATA1[30],DATA2[30],DATA3[30],SELECT,OUT[30],clk);
	MUX4x1 MUX31(DATA0[31],DATA1[31],DATA2[31],DATA3[31],SELECT,OUT[31],clk);
	MUX4x1 MUX32(DATA0[32],DATA1[32],DATA2[32],DATA3[32],SELECT,OUT[32],clk);
	MUX4x1 MUX33(DATA0[33],DATA1[33],DATA2[33],DATA3[33],SELECT,OUT[33],clk);
	MUX4x1 MUX34(DATA0[34],DATA1[34],DATA2[34],DATA3[34],SELECT,OUT[34],clk);
	MUX4x1 MUX35(DATA0[35],DATA1[35],DATA2[35],DATA3[35],SELECT,OUT[35],clk);
	MUX4x1 MUX36(DATA0[36],DATA1[36],DATA2[36],DATA3[36],SELECT,OUT[36],clk);
	MUX4x1 MUX37(DATA0[37],DATA1[37],DATA2[37],DATA3[37],SELECT,OUT[37],clk);
	MUX4x1 MUX38(DATA0[38],DATA1[38],DATA2[38],DATA3[38],SELECT,OUT[38],clk);
	MUX4x1 MUX39(DATA0[39],DATA1[39],DATA2[39],DATA3[39],SELECT,OUT[39],clk);
	MUX4x1 MUX40(DATA0[40],DATA1[40],DATA2[40],DATA3[40],SELECT,OUT[40],clk);
	MUX4x1 MUX41(DATA0[41],DATA1[41],DATA2[41],DATA3[41],SELECT,OUT[41],clk);
	MUX4x1 MUX42(DATA0[42],DATA1[42],DATA2[42],DATA3[42],SELECT,OUT[42],clk);
	MUX4x1 MUX43(DATA0[43],DATA1[43],DATA2[43],DATA3[43],SELECT,OUT[43],clk);
	MUX4x1 MUX44(DATA0[44],DATA1[44],DATA2[44],DATA3[44],SELECT,OUT[44],clk);
	MUX4x1 MUX45(DATA0[45],DATA1[45],DATA2[45],DATA3[45],SELECT,OUT[45],clk);
	MUX4x1 MUX46(DATA0[46],DATA1[46],DATA2[46],DATA3[46],SELECT,OUT[46],clk);
	MUX4x1 MUX47(DATA0[47],DATA1[47],DATA2[47],DATA3[47],SELECT,OUT[47],clk);
	MUX4x1 MUX48(DATA0[48],DATA1[48],DATA2[48],DATA3[48],SELECT,OUT[48],clk);
	MUX4x1 MUX49(DATA0[49],DATA1[49],DATA2[49],DATA3[49],SELECT,OUT[49],clk);
	MUX4x1 MUX50(DATA0[50],DATA1[50],DATA2[50],DATA3[50],SELECT,OUT[50],clk);
	MUX4x1 MUX51(DATA0[51],DATA1[51],DATA2[51],DATA3[51],SELECT,OUT[51],clk);
	MUX4x1 MUX52(DATA0[52],DATA1[52],DATA2[52],DATA3[52],SELECT,OUT[52],clk);
	MUX4x1 MUX53(DATA0[53],DATA1[53],DATA2[53],DATA3[53],SELECT,OUT[53],clk);
	MUX4x1 MUX54(DATA0[54],DATA1[54],DATA2[54],DATA3[54],SELECT,OUT[54],clk);
	MUX4x1 MUX55(DATA0[55],DATA1[55],DATA2[55],DATA3[55],SELECT,OUT[55],clk);
	MUX4x1 MUX56(DATA0[56],DATA1[56],DATA2[56],DATA3[56],SELECT,OUT[56],clk);
	MUX4x1 MUX57(DATA0[57],DATA1[57],DATA2[57],DATA3[57],SELECT,OUT[57],clk);
	MUX4x1 MUX58(DATA0[58],DATA1[58],DATA2[58],DATA3[58],SELECT,OUT[58],clk);
	MUX4x1 MUX59(DATA0[59],DATA1[59],DATA2[59],DATA3[59],SELECT,OUT[59],clk);
	MUX4x1 MUX60(DATA0[60],DATA1[60],DATA2[60],DATA3[60],SELECT,OUT[60],clk);
	MUX4x1 MUX61(DATA0[61],DATA1[61],DATA2[61],DATA3[61],SELECT,OUT[61],clk);
	MUX4x1 MUX62(DATA0[62],DATA1[62],DATA2[62],DATA3[62],SELECT,OUT[62],clk);
	MUX4x1 MUX63(DATA0[63],DATA1[63],DATA2[63],DATA3[63],SELECT,OUT[63],clk);
endmodule // MUX64bit_4x1

//2 stage Pipelined : 64 bit 4x1 MUX (For use in ALU)
//2 clock  cycles - input : clk 0; output : clk 2
module MUX64bit_16x1(DATA0,DATA1,DATA2,DATA3,DATA4,DATA5,DATA6,DATA7,DATA8,DATA9,DATA10,DATA11,DATA12,DATA13,DATA14,DATA15,SELECT,OUT,clk);

	input[63:0] DATA0,DATA1,DATA2,DATA3,DATA4,DATA5,DATA6,DATA7,DATA8,DATA9,DATA10,DATA11,DATA12,DATA13,DATA14,DATA15;
	input[3:0] SELECT;
	input clk;

	output[63:0] OUT;

	wire[63:0] LEVEL1_MUX0_OUT,LEVEL1_MUX1_OUT,LEVEL1_MUX2_OUT,LEVEL1_MUX3_OUT;
  	MUX64bit_4x1 level1_MUX0(DATA0,DATA1,DATA2,DATA3,SELECT[1:0],LEVEL1_MUX0_OUT,clk);
	MUX64bit_4x1 level1_MUX1(DATA4,DATA5,DATA6,DATA7,SELECT[1:0],LEVEL1_MUX1_OUT,clk);
	MUX64bit_4x1 level1_MUX2(DATA8,DATA9,DATA10,DATA11,SELECT[1:0],LEVEL1_MUX2_OUT,clk);
	MUX64bit_4x1 level1_MUX3(DATA12,DATA13,DATA14,DATA15,SELECT[1:0],LEVEL1_MUX3_OUT,clk);

	//Propogate MUX Outputs and select line values
	wire[63:0] LEVEL1_MUX0_FFOUT,LEVEL1_MUX1_FFOUT,LEVEL1_MUX2_FFOUT,LEVEL1_MUX3_FFOUT;
	DFlipFlop64 MUX0_outFF(LEVEL1_MUX0_OUT,clk,LEVEL1_MUX0_FFOUT);
	DFlipFlop64 MUX1_outFF(LEVEL1_MUX1_OUT,clk,LEVEL1_MUX1_FFOUT);
	DFlipFlop64 MUX2_outFF(LEVEL1_MUX2_OUT,clk,LEVEL1_MUX2_FFOUT);
	DFlipFlop64 MUX3_outFF(LEVEL1_MUX3_OUT,clk,LEVEL1_MUX3_FFOUT);

	wire[1:0] LEVEL1_SELECT_FFOUT;
	DFlipFlop2 level1_SELECT_FF(SELECT[3:2],clk,LEVEL1_SELECT_FFOUT);

	MUX64bit_4x1 level2_MUX(LEVEL1_MUX0_FFOUT,LEVEL1_MUX1_FFOUT,LEVEL1_MUX2_FFOUT,LEVEL1_MUX3_FFOUT,LEVEL1_SELECT_FFOUT,OUT,clk);

endmodule // MUX64bit_16x1

`endif
