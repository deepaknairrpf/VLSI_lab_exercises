//header guards
`ifndef _memory_vh_
`define _memory_vh_


`include "decoders.v"
`include "tristate.v"
`include "DFFwithEnable.v"

//Should we able to read and write at same time?
module memory256x32bit(cs,rd_wr,ADDRESS,DATAIN,DATAOUT,clk);

	//inputs: CHIP SELECT, read/~write 
	input cs,rd_wr,clk;
	input[7:0] ADDRESS;
	input[31:0] DATAIN;

	output[31:0] DATAOUT;

	wire[255:0] DECODER_OUT;

	wire[31:0] DFF_OUT[0:255];

	decoder8x256 decoder(cs,ADDRESS,DECODER_OUT);

  //DFF32bitEnable DFF0(DATAIN,clk,DFF_OUT[0],DECODER_OUT[0]&~rd_wr);
  	//WRITING TO MEMORY
	DFF32bitEnable DFF0(DATAIN,clk,DFF_OUT[0],DECODER_OUT[0]&~rd_wr);
	DFF32bitEnable DFF1(DATAIN,clk,DFF_OUT[1],DECODER_OUT[1]&~rd_wr);
	DFF32bitEnable DFF2(DATAIN,clk,DFF_OUT[2],DECODER_OUT[2]&~rd_wr);
	DFF32bitEnable DFF3(DATAIN,clk,DFF_OUT[3],DECODER_OUT[3]&~rd_wr);
	DFF32bitEnable DFF4(DATAIN,clk,DFF_OUT[4],DECODER_OUT[4]&~rd_wr);
	DFF32bitEnable DFF5(DATAIN,clk,DFF_OUT[5],DECODER_OUT[5]&~rd_wr);
	DFF32bitEnable DFF6(DATAIN,clk,DFF_OUT[6],DECODER_OUT[6]&~rd_wr);
	DFF32bitEnable DFF7(DATAIN,clk,DFF_OUT[7],DECODER_OUT[7]&~rd_wr);
	DFF32bitEnable DFF8(DATAIN,clk,DFF_OUT[8],DECODER_OUT[8]&~rd_wr);
	DFF32bitEnable DFF9(DATAIN,clk,DFF_OUT[9],DECODER_OUT[9]&~rd_wr);
	DFF32bitEnable DFF10(DATAIN,clk,DFF_OUT[10],DECODER_OUT[10]&~rd_wr);
	DFF32bitEnable DFF11(DATAIN,clk,DFF_OUT[11],DECODER_OUT[11]&~rd_wr);
	DFF32bitEnable DFF12(DATAIN,clk,DFF_OUT[12],DECODER_OUT[12]&~rd_wr);
	DFF32bitEnable DFF13(DATAIN,clk,DFF_OUT[13],DECODER_OUT[13]&~rd_wr);
	DFF32bitEnable DFF14(DATAIN,clk,DFF_OUT[14],DECODER_OUT[14]&~rd_wr);
	DFF32bitEnable DFF15(DATAIN,clk,DFF_OUT[15],DECODER_OUT[15]&~rd_wr);
	DFF32bitEnable DFF16(DATAIN,clk,DFF_OUT[16],DECODER_OUT[16]&~rd_wr);
	DFF32bitEnable DFF17(DATAIN,clk,DFF_OUT[17],DECODER_OUT[17]&~rd_wr);
	DFF32bitEnable DFF18(DATAIN,clk,DFF_OUT[18],DECODER_OUT[18]&~rd_wr);
	DFF32bitEnable DFF19(DATAIN,clk,DFF_OUT[19],DECODER_OUT[19]&~rd_wr);
	DFF32bitEnable DFF20(DATAIN,clk,DFF_OUT[20],DECODER_OUT[20]&~rd_wr);
	DFF32bitEnable DFF21(DATAIN,clk,DFF_OUT[21],DECODER_OUT[21]&~rd_wr);
	DFF32bitEnable DFF22(DATAIN,clk,DFF_OUT[22],DECODER_OUT[22]&~rd_wr);
	DFF32bitEnable DFF23(DATAIN,clk,DFF_OUT[23],DECODER_OUT[23]&~rd_wr);
	DFF32bitEnable DFF24(DATAIN,clk,DFF_OUT[24],DECODER_OUT[24]&~rd_wr);
	DFF32bitEnable DFF25(DATAIN,clk,DFF_OUT[25],DECODER_OUT[25]&~rd_wr);
	DFF32bitEnable DFF26(DATAIN,clk,DFF_OUT[26],DECODER_OUT[26]&~rd_wr);
	DFF32bitEnable DFF27(DATAIN,clk,DFF_OUT[27],DECODER_OUT[27]&~rd_wr);
	DFF32bitEnable DFF28(DATAIN,clk,DFF_OUT[28],DECODER_OUT[28]&~rd_wr);
	DFF32bitEnable DFF29(DATAIN,clk,DFF_OUT[29],DECODER_OUT[29]&~rd_wr);
	DFF32bitEnable DFF30(DATAIN,clk,DFF_OUT[30],DECODER_OUT[30]&~rd_wr);
	DFF32bitEnable DFF31(DATAIN,clk,DFF_OUT[31],DECODER_OUT[31]&~rd_wr);
	DFF32bitEnable DFF32(DATAIN,clk,DFF_OUT[32],DECODER_OUT[32]&~rd_wr);
	DFF32bitEnable DFF33(DATAIN,clk,DFF_OUT[33],DECODER_OUT[33]&~rd_wr);
	DFF32bitEnable DFF34(DATAIN,clk,DFF_OUT[34],DECODER_OUT[34]&~rd_wr);
	DFF32bitEnable DFF35(DATAIN,clk,DFF_OUT[35],DECODER_OUT[35]&~rd_wr);
	DFF32bitEnable DFF36(DATAIN,clk,DFF_OUT[36],DECODER_OUT[36]&~rd_wr);
	DFF32bitEnable DFF37(DATAIN,clk,DFF_OUT[37],DECODER_OUT[37]&~rd_wr);
	DFF32bitEnable DFF38(DATAIN,clk,DFF_OUT[38],DECODER_OUT[38]&~rd_wr);
	DFF32bitEnable DFF39(DATAIN,clk,DFF_OUT[39],DECODER_OUT[39]&~rd_wr);
	DFF32bitEnable DFF40(DATAIN,clk,DFF_OUT[40],DECODER_OUT[40]&~rd_wr);
	DFF32bitEnable DFF41(DATAIN,clk,DFF_OUT[41],DECODER_OUT[41]&~rd_wr);
	DFF32bitEnable DFF42(DATAIN,clk,DFF_OUT[42],DECODER_OUT[42]&~rd_wr);
	DFF32bitEnable DFF43(DATAIN,clk,DFF_OUT[43],DECODER_OUT[43]&~rd_wr);
	DFF32bitEnable DFF44(DATAIN,clk,DFF_OUT[44],DECODER_OUT[44]&~rd_wr);
	DFF32bitEnable DFF45(DATAIN,clk,DFF_OUT[45],DECODER_OUT[45]&~rd_wr);
	DFF32bitEnable DFF46(DATAIN,clk,DFF_OUT[46],DECODER_OUT[46]&~rd_wr);
	DFF32bitEnable DFF47(DATAIN,clk,DFF_OUT[47],DECODER_OUT[47]&~rd_wr);
	DFF32bitEnable DFF48(DATAIN,clk,DFF_OUT[48],DECODER_OUT[48]&~rd_wr);
	DFF32bitEnable DFF49(DATAIN,clk,DFF_OUT[49],DECODER_OUT[49]&~rd_wr);
	DFF32bitEnable DFF50(DATAIN,clk,DFF_OUT[50],DECODER_OUT[50]&~rd_wr);
	DFF32bitEnable DFF51(DATAIN,clk,DFF_OUT[51],DECODER_OUT[51]&~rd_wr);
	DFF32bitEnable DFF52(DATAIN,clk,DFF_OUT[52],DECODER_OUT[52]&~rd_wr);
	DFF32bitEnable DFF53(DATAIN,clk,DFF_OUT[53],DECODER_OUT[53]&~rd_wr);
	DFF32bitEnable DFF54(DATAIN,clk,DFF_OUT[54],DECODER_OUT[54]&~rd_wr);
	DFF32bitEnable DFF55(DATAIN,clk,DFF_OUT[55],DECODER_OUT[55]&~rd_wr);
	DFF32bitEnable DFF56(DATAIN,clk,DFF_OUT[56],DECODER_OUT[56]&~rd_wr);
	DFF32bitEnable DFF57(DATAIN,clk,DFF_OUT[57],DECODER_OUT[57]&~rd_wr);
	DFF32bitEnable DFF58(DATAIN,clk,DFF_OUT[58],DECODER_OUT[58]&~rd_wr);
	DFF32bitEnable DFF59(DATAIN,clk,DFF_OUT[59],DECODER_OUT[59]&~rd_wr);
	DFF32bitEnable DFF60(DATAIN,clk,DFF_OUT[60],DECODER_OUT[60]&~rd_wr);
	DFF32bitEnable DFF61(DATAIN,clk,DFF_OUT[61],DECODER_OUT[61]&~rd_wr);
	DFF32bitEnable DFF62(DATAIN,clk,DFF_OUT[62],DECODER_OUT[62]&~rd_wr);
	DFF32bitEnable DFF63(DATAIN,clk,DFF_OUT[63],DECODER_OUT[63]&~rd_wr);
	DFF32bitEnable DFF64(DATAIN,clk,DFF_OUT[64],DECODER_OUT[64]&~rd_wr);
	DFF32bitEnable DFF65(DATAIN,clk,DFF_OUT[65],DECODER_OUT[65]&~rd_wr);
	DFF32bitEnable DFF66(DATAIN,clk,DFF_OUT[66],DECODER_OUT[66]&~rd_wr);
	DFF32bitEnable DFF67(DATAIN,clk,DFF_OUT[67],DECODER_OUT[67]&~rd_wr);
	DFF32bitEnable DFF68(DATAIN,clk,DFF_OUT[68],DECODER_OUT[68]&~rd_wr);
	DFF32bitEnable DFF69(DATAIN,clk,DFF_OUT[69],DECODER_OUT[69]&~rd_wr);
	DFF32bitEnable DFF70(DATAIN,clk,DFF_OUT[70],DECODER_OUT[70]&~rd_wr);
	DFF32bitEnable DFF71(DATAIN,clk,DFF_OUT[71],DECODER_OUT[71]&~rd_wr);
	DFF32bitEnable DFF72(DATAIN,clk,DFF_OUT[72],DECODER_OUT[72]&~rd_wr);
	DFF32bitEnable DFF73(DATAIN,clk,DFF_OUT[73],DECODER_OUT[73]&~rd_wr);
	DFF32bitEnable DFF74(DATAIN,clk,DFF_OUT[74],DECODER_OUT[74]&~rd_wr);
	DFF32bitEnable DFF75(DATAIN,clk,DFF_OUT[75],DECODER_OUT[75]&~rd_wr);
	DFF32bitEnable DFF76(DATAIN,clk,DFF_OUT[76],DECODER_OUT[76]&~rd_wr);
	DFF32bitEnable DFF77(DATAIN,clk,DFF_OUT[77],DECODER_OUT[77]&~rd_wr);
	DFF32bitEnable DFF78(DATAIN,clk,DFF_OUT[78],DECODER_OUT[78]&~rd_wr);
	DFF32bitEnable DFF79(DATAIN,clk,DFF_OUT[79],DECODER_OUT[79]&~rd_wr);
	DFF32bitEnable DFF80(DATAIN,clk,DFF_OUT[80],DECODER_OUT[80]&~rd_wr);
	DFF32bitEnable DFF81(DATAIN,clk,DFF_OUT[81],DECODER_OUT[81]&~rd_wr);
	DFF32bitEnable DFF82(DATAIN,clk,DFF_OUT[82],DECODER_OUT[82]&~rd_wr);
	DFF32bitEnable DFF83(DATAIN,clk,DFF_OUT[83],DECODER_OUT[83]&~rd_wr);
	DFF32bitEnable DFF84(DATAIN,clk,DFF_OUT[84],DECODER_OUT[84]&~rd_wr);
	DFF32bitEnable DFF85(DATAIN,clk,DFF_OUT[85],DECODER_OUT[85]&~rd_wr);
	DFF32bitEnable DFF86(DATAIN,clk,DFF_OUT[86],DECODER_OUT[86]&~rd_wr);
	DFF32bitEnable DFF87(DATAIN,clk,DFF_OUT[87],DECODER_OUT[87]&~rd_wr);
	DFF32bitEnable DFF88(DATAIN,clk,DFF_OUT[88],DECODER_OUT[88]&~rd_wr);
	DFF32bitEnable DFF89(DATAIN,clk,DFF_OUT[89],DECODER_OUT[89]&~rd_wr);
	DFF32bitEnable DFF90(DATAIN,clk,DFF_OUT[90],DECODER_OUT[90]&~rd_wr);
	DFF32bitEnable DFF91(DATAIN,clk,DFF_OUT[91],DECODER_OUT[91]&~rd_wr);
	DFF32bitEnable DFF92(DATAIN,clk,DFF_OUT[92],DECODER_OUT[92]&~rd_wr);
	DFF32bitEnable DFF93(DATAIN,clk,DFF_OUT[93],DECODER_OUT[93]&~rd_wr);
	DFF32bitEnable DFF94(DATAIN,clk,DFF_OUT[94],DECODER_OUT[94]&~rd_wr);
	DFF32bitEnable DFF95(DATAIN,clk,DFF_OUT[95],DECODER_OUT[95]&~rd_wr);
	DFF32bitEnable DFF96(DATAIN,clk,DFF_OUT[96],DECODER_OUT[96]&~rd_wr);
	DFF32bitEnable DFF97(DATAIN,clk,DFF_OUT[97],DECODER_OUT[97]&~rd_wr);
	DFF32bitEnable DFF98(DATAIN,clk,DFF_OUT[98],DECODER_OUT[98]&~rd_wr);
	DFF32bitEnable DFF99(DATAIN,clk,DFF_OUT[99],DECODER_OUT[99]&~rd_wr);
	DFF32bitEnable DFF100(DATAIN,clk,DFF_OUT[100],DECODER_OUT[100]&~rd_wr);
	DFF32bitEnable DFF101(DATAIN,clk,DFF_OUT[101],DECODER_OUT[101]&~rd_wr);
	DFF32bitEnable DFF102(DATAIN,clk,DFF_OUT[102],DECODER_OUT[102]&~rd_wr);
	DFF32bitEnable DFF103(DATAIN,clk,DFF_OUT[103],DECODER_OUT[103]&~rd_wr);
	DFF32bitEnable DFF104(DATAIN,clk,DFF_OUT[104],DECODER_OUT[104]&~rd_wr);
	DFF32bitEnable DFF105(DATAIN,clk,DFF_OUT[105],DECODER_OUT[105]&~rd_wr);
	DFF32bitEnable DFF106(DATAIN,clk,DFF_OUT[106],DECODER_OUT[106]&~rd_wr);
	DFF32bitEnable DFF107(DATAIN,clk,DFF_OUT[107],DECODER_OUT[107]&~rd_wr);
	DFF32bitEnable DFF108(DATAIN,clk,DFF_OUT[108],DECODER_OUT[108]&~rd_wr);
	DFF32bitEnable DFF109(DATAIN,clk,DFF_OUT[109],DECODER_OUT[109]&~rd_wr);
	DFF32bitEnable DFF110(DATAIN,clk,DFF_OUT[110],DECODER_OUT[110]&~rd_wr);
	DFF32bitEnable DFF111(DATAIN,clk,DFF_OUT[111],DECODER_OUT[111]&~rd_wr);
	DFF32bitEnable DFF112(DATAIN,clk,DFF_OUT[112],DECODER_OUT[112]&~rd_wr);
	DFF32bitEnable DFF113(DATAIN,clk,DFF_OUT[113],DECODER_OUT[113]&~rd_wr);
	DFF32bitEnable DFF114(DATAIN,clk,DFF_OUT[114],DECODER_OUT[114]&~rd_wr);
	DFF32bitEnable DFF115(DATAIN,clk,DFF_OUT[115],DECODER_OUT[115]&~rd_wr);
	DFF32bitEnable DFF116(DATAIN,clk,DFF_OUT[116],DECODER_OUT[116]&~rd_wr);
	DFF32bitEnable DFF117(DATAIN,clk,DFF_OUT[117],DECODER_OUT[117]&~rd_wr);
	DFF32bitEnable DFF118(DATAIN,clk,DFF_OUT[118],DECODER_OUT[118]&~rd_wr);
	DFF32bitEnable DFF119(DATAIN,clk,DFF_OUT[119],DECODER_OUT[119]&~rd_wr);
	DFF32bitEnable DFF120(DATAIN,clk,DFF_OUT[120],DECODER_OUT[120]&~rd_wr);
	DFF32bitEnable DFF121(DATAIN,clk,DFF_OUT[121],DECODER_OUT[121]&~rd_wr);
	DFF32bitEnable DFF122(DATAIN,clk,DFF_OUT[122],DECODER_OUT[122]&~rd_wr);
	DFF32bitEnable DFF123(DATAIN,clk,DFF_OUT[123],DECODER_OUT[123]&~rd_wr);
	DFF32bitEnable DFF124(DATAIN,clk,DFF_OUT[124],DECODER_OUT[124]&~rd_wr);
	DFF32bitEnable DFF125(DATAIN,clk,DFF_OUT[125],DECODER_OUT[125]&~rd_wr);
	DFF32bitEnable DFF126(DATAIN,clk,DFF_OUT[126],DECODER_OUT[126]&~rd_wr);
	DFF32bitEnable DFF127(DATAIN,clk,DFF_OUT[127],DECODER_OUT[127]&~rd_wr);
	DFF32bitEnable DFF128(DATAIN,clk,DFF_OUT[128],DECODER_OUT[128]&~rd_wr);
	DFF32bitEnable DFF129(DATAIN,clk,DFF_OUT[129],DECODER_OUT[129]&~rd_wr);
	DFF32bitEnable DFF130(DATAIN,clk,DFF_OUT[130],DECODER_OUT[130]&~rd_wr);
	DFF32bitEnable DFF131(DATAIN,clk,DFF_OUT[131],DECODER_OUT[131]&~rd_wr);
	DFF32bitEnable DFF132(DATAIN,clk,DFF_OUT[132],DECODER_OUT[132]&~rd_wr);
	DFF32bitEnable DFF133(DATAIN,clk,DFF_OUT[133],DECODER_OUT[133]&~rd_wr);
	DFF32bitEnable DFF134(DATAIN,clk,DFF_OUT[134],DECODER_OUT[134]&~rd_wr);
	DFF32bitEnable DFF135(DATAIN,clk,DFF_OUT[135],DECODER_OUT[135]&~rd_wr);
	DFF32bitEnable DFF136(DATAIN,clk,DFF_OUT[136],DECODER_OUT[136]&~rd_wr);
	DFF32bitEnable DFF137(DATAIN,clk,DFF_OUT[137],DECODER_OUT[137]&~rd_wr);
	DFF32bitEnable DFF138(DATAIN,clk,DFF_OUT[138],DECODER_OUT[138]&~rd_wr);
	DFF32bitEnable DFF139(DATAIN,clk,DFF_OUT[139],DECODER_OUT[139]&~rd_wr);
	DFF32bitEnable DFF140(DATAIN,clk,DFF_OUT[140],DECODER_OUT[140]&~rd_wr);
	DFF32bitEnable DFF141(DATAIN,clk,DFF_OUT[141],DECODER_OUT[141]&~rd_wr);
	DFF32bitEnable DFF142(DATAIN,clk,DFF_OUT[142],DECODER_OUT[142]&~rd_wr);
	DFF32bitEnable DFF143(DATAIN,clk,DFF_OUT[143],DECODER_OUT[143]&~rd_wr);
	DFF32bitEnable DFF144(DATAIN,clk,DFF_OUT[144],DECODER_OUT[144]&~rd_wr);
	DFF32bitEnable DFF145(DATAIN,clk,DFF_OUT[145],DECODER_OUT[145]&~rd_wr);
	DFF32bitEnable DFF146(DATAIN,clk,DFF_OUT[146],DECODER_OUT[146]&~rd_wr);
	DFF32bitEnable DFF147(DATAIN,clk,DFF_OUT[147],DECODER_OUT[147]&~rd_wr);
	DFF32bitEnable DFF148(DATAIN,clk,DFF_OUT[148],DECODER_OUT[148]&~rd_wr);
	DFF32bitEnable DFF149(DATAIN,clk,DFF_OUT[149],DECODER_OUT[149]&~rd_wr);
	DFF32bitEnable DFF150(DATAIN,clk,DFF_OUT[150],DECODER_OUT[150]&~rd_wr);
	DFF32bitEnable DFF151(DATAIN,clk,DFF_OUT[151],DECODER_OUT[151]&~rd_wr);
	DFF32bitEnable DFF152(DATAIN,clk,DFF_OUT[152],DECODER_OUT[152]&~rd_wr);
	DFF32bitEnable DFF153(DATAIN,clk,DFF_OUT[153],DECODER_OUT[153]&~rd_wr);
	DFF32bitEnable DFF154(DATAIN,clk,DFF_OUT[154],DECODER_OUT[154]&~rd_wr);
	DFF32bitEnable DFF155(DATAIN,clk,DFF_OUT[155],DECODER_OUT[155]&~rd_wr);
	DFF32bitEnable DFF156(DATAIN,clk,DFF_OUT[156],DECODER_OUT[156]&~rd_wr);
	DFF32bitEnable DFF157(DATAIN,clk,DFF_OUT[157],DECODER_OUT[157]&~rd_wr);
	DFF32bitEnable DFF158(DATAIN,clk,DFF_OUT[158],DECODER_OUT[158]&~rd_wr);
	DFF32bitEnable DFF159(DATAIN,clk,DFF_OUT[159],DECODER_OUT[159]&~rd_wr);
	DFF32bitEnable DFF160(DATAIN,clk,DFF_OUT[160],DECODER_OUT[160]&~rd_wr);
	DFF32bitEnable DFF161(DATAIN,clk,DFF_OUT[161],DECODER_OUT[161]&~rd_wr);
	DFF32bitEnable DFF162(DATAIN,clk,DFF_OUT[162],DECODER_OUT[162]&~rd_wr);
	DFF32bitEnable DFF163(DATAIN,clk,DFF_OUT[163],DECODER_OUT[163]&~rd_wr);
	DFF32bitEnable DFF164(DATAIN,clk,DFF_OUT[164],DECODER_OUT[164]&~rd_wr);
	DFF32bitEnable DFF165(DATAIN,clk,DFF_OUT[165],DECODER_OUT[165]&~rd_wr);
	DFF32bitEnable DFF166(DATAIN,clk,DFF_OUT[166],DECODER_OUT[166]&~rd_wr);
	DFF32bitEnable DFF167(DATAIN,clk,DFF_OUT[167],DECODER_OUT[167]&~rd_wr);
	DFF32bitEnable DFF168(DATAIN,clk,DFF_OUT[168],DECODER_OUT[168]&~rd_wr);
	DFF32bitEnable DFF169(DATAIN,clk,DFF_OUT[169],DECODER_OUT[169]&~rd_wr);
	DFF32bitEnable DFF170(DATAIN,clk,DFF_OUT[170],DECODER_OUT[170]&~rd_wr);
	DFF32bitEnable DFF171(DATAIN,clk,DFF_OUT[171],DECODER_OUT[171]&~rd_wr);
	DFF32bitEnable DFF172(DATAIN,clk,DFF_OUT[172],DECODER_OUT[172]&~rd_wr);
	DFF32bitEnable DFF173(DATAIN,clk,DFF_OUT[173],DECODER_OUT[173]&~rd_wr);
	DFF32bitEnable DFF174(DATAIN,clk,DFF_OUT[174],DECODER_OUT[174]&~rd_wr);
	DFF32bitEnable DFF175(DATAIN,clk,DFF_OUT[175],DECODER_OUT[175]&~rd_wr);
	DFF32bitEnable DFF176(DATAIN,clk,DFF_OUT[176],DECODER_OUT[176]&~rd_wr);
	DFF32bitEnable DFF177(DATAIN,clk,DFF_OUT[177],DECODER_OUT[177]&~rd_wr);
	DFF32bitEnable DFF178(DATAIN,clk,DFF_OUT[178],DECODER_OUT[178]&~rd_wr);
	DFF32bitEnable DFF179(DATAIN,clk,DFF_OUT[179],DECODER_OUT[179]&~rd_wr);
	DFF32bitEnable DFF180(DATAIN,clk,DFF_OUT[180],DECODER_OUT[180]&~rd_wr);
	DFF32bitEnable DFF181(DATAIN,clk,DFF_OUT[181],DECODER_OUT[181]&~rd_wr);
	DFF32bitEnable DFF182(DATAIN,clk,DFF_OUT[182],DECODER_OUT[182]&~rd_wr);
	DFF32bitEnable DFF183(DATAIN,clk,DFF_OUT[183],DECODER_OUT[183]&~rd_wr);
	DFF32bitEnable DFF184(DATAIN,clk,DFF_OUT[184],DECODER_OUT[184]&~rd_wr);
	DFF32bitEnable DFF185(DATAIN,clk,DFF_OUT[185],DECODER_OUT[185]&~rd_wr);
	DFF32bitEnable DFF186(DATAIN,clk,DFF_OUT[186],DECODER_OUT[186]&~rd_wr);
	DFF32bitEnable DFF187(DATAIN,clk,DFF_OUT[187],DECODER_OUT[187]&~rd_wr);
	DFF32bitEnable DFF188(DATAIN,clk,DFF_OUT[188],DECODER_OUT[188]&~rd_wr);
	DFF32bitEnable DFF189(DATAIN,clk,DFF_OUT[189],DECODER_OUT[189]&~rd_wr);
	DFF32bitEnable DFF190(DATAIN,clk,DFF_OUT[190],DECODER_OUT[190]&~rd_wr);
	DFF32bitEnable DFF191(DATAIN,clk,DFF_OUT[191],DECODER_OUT[191]&~rd_wr);
	DFF32bitEnable DFF192(DATAIN,clk,DFF_OUT[192],DECODER_OUT[192]&~rd_wr);
	DFF32bitEnable DFF193(DATAIN,clk,DFF_OUT[193],DECODER_OUT[193]&~rd_wr);
	DFF32bitEnable DFF194(DATAIN,clk,DFF_OUT[194],DECODER_OUT[194]&~rd_wr);
	DFF32bitEnable DFF195(DATAIN,clk,DFF_OUT[195],DECODER_OUT[195]&~rd_wr);
	DFF32bitEnable DFF196(DATAIN,clk,DFF_OUT[196],DECODER_OUT[196]&~rd_wr);
	DFF32bitEnable DFF197(DATAIN,clk,DFF_OUT[197],DECODER_OUT[197]&~rd_wr);
	DFF32bitEnable DFF198(DATAIN,clk,DFF_OUT[198],DECODER_OUT[198]&~rd_wr);
	DFF32bitEnable DFF199(DATAIN,clk,DFF_OUT[199],DECODER_OUT[199]&~rd_wr);
	DFF32bitEnable DFF200(DATAIN,clk,DFF_OUT[200],DECODER_OUT[200]&~rd_wr);
	DFF32bitEnable DFF201(DATAIN,clk,DFF_OUT[201],DECODER_OUT[201]&~rd_wr);
	DFF32bitEnable DFF202(DATAIN,clk,DFF_OUT[202],DECODER_OUT[202]&~rd_wr);
	DFF32bitEnable DFF203(DATAIN,clk,DFF_OUT[203],DECODER_OUT[203]&~rd_wr);
	DFF32bitEnable DFF204(DATAIN,clk,DFF_OUT[204],DECODER_OUT[204]&~rd_wr);
	DFF32bitEnable DFF205(DATAIN,clk,DFF_OUT[205],DECODER_OUT[205]&~rd_wr);
	DFF32bitEnable DFF206(DATAIN,clk,DFF_OUT[206],DECODER_OUT[206]&~rd_wr);
	DFF32bitEnable DFF207(DATAIN,clk,DFF_OUT[207],DECODER_OUT[207]&~rd_wr);
	DFF32bitEnable DFF208(DATAIN,clk,DFF_OUT[208],DECODER_OUT[208]&~rd_wr);
	DFF32bitEnable DFF209(DATAIN,clk,DFF_OUT[209],DECODER_OUT[209]&~rd_wr);
	DFF32bitEnable DFF210(DATAIN,clk,DFF_OUT[210],DECODER_OUT[210]&~rd_wr);
	DFF32bitEnable DFF211(DATAIN,clk,DFF_OUT[211],DECODER_OUT[211]&~rd_wr);
	DFF32bitEnable DFF212(DATAIN,clk,DFF_OUT[212],DECODER_OUT[212]&~rd_wr);
	DFF32bitEnable DFF213(DATAIN,clk,DFF_OUT[213],DECODER_OUT[213]&~rd_wr);
	DFF32bitEnable DFF214(DATAIN,clk,DFF_OUT[214],DECODER_OUT[214]&~rd_wr);
	DFF32bitEnable DFF215(DATAIN,clk,DFF_OUT[215],DECODER_OUT[215]&~rd_wr);
	DFF32bitEnable DFF216(DATAIN,clk,DFF_OUT[216],DECODER_OUT[216]&~rd_wr);
	DFF32bitEnable DFF217(DATAIN,clk,DFF_OUT[217],DECODER_OUT[217]&~rd_wr);
	DFF32bitEnable DFF218(DATAIN,clk,DFF_OUT[218],DECODER_OUT[218]&~rd_wr);
	DFF32bitEnable DFF219(DATAIN,clk,DFF_OUT[219],DECODER_OUT[219]&~rd_wr);
	DFF32bitEnable DFF220(DATAIN,clk,DFF_OUT[220],DECODER_OUT[220]&~rd_wr);
	DFF32bitEnable DFF221(DATAIN,clk,DFF_OUT[221],DECODER_OUT[221]&~rd_wr);
	DFF32bitEnable DFF222(DATAIN,clk,DFF_OUT[222],DECODER_OUT[222]&~rd_wr);
	DFF32bitEnable DFF223(DATAIN,clk,DFF_OUT[223],DECODER_OUT[223]&~rd_wr);
	DFF32bitEnable DFF224(DATAIN,clk,DFF_OUT[224],DECODER_OUT[224]&~rd_wr);
	DFF32bitEnable DFF225(DATAIN,clk,DFF_OUT[225],DECODER_OUT[225]&~rd_wr);
	DFF32bitEnable DFF226(DATAIN,clk,DFF_OUT[226],DECODER_OUT[226]&~rd_wr);
	DFF32bitEnable DFF227(DATAIN,clk,DFF_OUT[227],DECODER_OUT[227]&~rd_wr);
	DFF32bitEnable DFF228(DATAIN,clk,DFF_OUT[228],DECODER_OUT[228]&~rd_wr);
	DFF32bitEnable DFF229(DATAIN,clk,DFF_OUT[229],DECODER_OUT[229]&~rd_wr);
	DFF32bitEnable DFF230(DATAIN,clk,DFF_OUT[230],DECODER_OUT[230]&~rd_wr);
	DFF32bitEnable DFF231(DATAIN,clk,DFF_OUT[231],DECODER_OUT[231]&~rd_wr);
	DFF32bitEnable DFF232(DATAIN,clk,DFF_OUT[232],DECODER_OUT[232]&~rd_wr);
	DFF32bitEnable DFF233(DATAIN,clk,DFF_OUT[233],DECODER_OUT[233]&~rd_wr);
	DFF32bitEnable DFF234(DATAIN,clk,DFF_OUT[234],DECODER_OUT[234]&~rd_wr);
	DFF32bitEnable DFF235(DATAIN,clk,DFF_OUT[235],DECODER_OUT[235]&~rd_wr);
	DFF32bitEnable DFF236(DATAIN,clk,DFF_OUT[236],DECODER_OUT[236]&~rd_wr);
	DFF32bitEnable DFF237(DATAIN,clk,DFF_OUT[237],DECODER_OUT[237]&~rd_wr);
	DFF32bitEnable DFF238(DATAIN,clk,DFF_OUT[238],DECODER_OUT[238]&~rd_wr);
	DFF32bitEnable DFF239(DATAIN,clk,DFF_OUT[239],DECODER_OUT[239]&~rd_wr);
	DFF32bitEnable DFF240(DATAIN,clk,DFF_OUT[240],DECODER_OUT[240]&~rd_wr);
	DFF32bitEnable DFF241(DATAIN,clk,DFF_OUT[241],DECODER_OUT[241]&~rd_wr);
	DFF32bitEnable DFF242(DATAIN,clk,DFF_OUT[242],DECODER_OUT[242]&~rd_wr);
	DFF32bitEnable DFF243(DATAIN,clk,DFF_OUT[243],DECODER_OUT[243]&~rd_wr);
	DFF32bitEnable DFF244(DATAIN,clk,DFF_OUT[244],DECODER_OUT[244]&~rd_wr);
	DFF32bitEnable DFF245(DATAIN,clk,DFF_OUT[245],DECODER_OUT[245]&~rd_wr);
	DFF32bitEnable DFF246(DATAIN,clk,DFF_OUT[246],DECODER_OUT[246]&~rd_wr);
	DFF32bitEnable DFF247(DATAIN,clk,DFF_OUT[247],DECODER_OUT[247]&~rd_wr);
	DFF32bitEnable DFF248(DATAIN,clk,DFF_OUT[248],DECODER_OUT[248]&~rd_wr);
	DFF32bitEnable DFF249(DATAIN,clk,DFF_OUT[249],DECODER_OUT[249]&~rd_wr);
	DFF32bitEnable DFF250(DATAIN,clk,DFF_OUT[250],DECODER_OUT[250]&~rd_wr);
	DFF32bitEnable DFF251(DATAIN,clk,DFF_OUT[251],DECODER_OUT[251]&~rd_wr);
	DFF32bitEnable DFF252(DATAIN,clk,DFF_OUT[252],DECODER_OUT[252]&~rd_wr);
	DFF32bitEnable DFF253(DATAIN,clk,DFF_OUT[253],DECODER_OUT[253]&~rd_wr);
	DFF32bitEnable DFF254(DATAIN,clk,DFF_OUT[254],DECODER_OUT[254]&~rd_wr);
	DFF32bitEnable DFF255(DATAIN,clk,DFF_OUT[255],DECODER_OUT[255]&~rd_wr);

	//READING FROM MEMORY
    //tristate32bit TSB0(DFF_OUT[0],DECODER_OUT[0]&rd_wr,DATAOUT);

	tristate32bit TSB0(DFF_OUT[0],DECODER_OUT[0]&rd_wr,DATAOUT);
	tristate32bit TSB1(DFF_OUT[1],DECODER_OUT[1]&rd_wr,DATAOUT);
	tristate32bit TSB2(DFF_OUT[2],DECODER_OUT[2]&rd_wr,DATAOUT);
	tristate32bit TSB3(DFF_OUT[3],DECODER_OUT[3]&rd_wr,DATAOUT);
	tristate32bit TSB4(DFF_OUT[4],DECODER_OUT[4]&rd_wr,DATAOUT);
	tristate32bit TSB5(DFF_OUT[5],DECODER_OUT[5]&rd_wr,DATAOUT);
	tristate32bit TSB6(DFF_OUT[6],DECODER_OUT[6]&rd_wr,DATAOUT);
	tristate32bit TSB7(DFF_OUT[7],DECODER_OUT[7]&rd_wr,DATAOUT);
	tristate32bit TSB8(DFF_OUT[8],DECODER_OUT[8]&rd_wr,DATAOUT);
	tristate32bit TSB9(DFF_OUT[9],DECODER_OUT[9]&rd_wr,DATAOUT);
	tristate32bit TSB10(DFF_OUT[10],DECODER_OUT[10]&rd_wr,DATAOUT);
	tristate32bit TSB11(DFF_OUT[11],DECODER_OUT[11]&rd_wr,DATAOUT);
	tristate32bit TSB12(DFF_OUT[12],DECODER_OUT[12]&rd_wr,DATAOUT);
	tristate32bit TSB13(DFF_OUT[13],DECODER_OUT[13]&rd_wr,DATAOUT);
	tristate32bit TSB14(DFF_OUT[14],DECODER_OUT[14]&rd_wr,DATAOUT);
	tristate32bit TSB15(DFF_OUT[15],DECODER_OUT[15]&rd_wr,DATAOUT);
	tristate32bit TSB16(DFF_OUT[16],DECODER_OUT[16]&rd_wr,DATAOUT);
	tristate32bit TSB17(DFF_OUT[17],DECODER_OUT[17]&rd_wr,DATAOUT);
	tristate32bit TSB18(DFF_OUT[18],DECODER_OUT[18]&rd_wr,DATAOUT);
	tristate32bit TSB19(DFF_OUT[19],DECODER_OUT[19]&rd_wr,DATAOUT);
	tristate32bit TSB20(DFF_OUT[20],DECODER_OUT[20]&rd_wr,DATAOUT);
	tristate32bit TSB21(DFF_OUT[21],DECODER_OUT[21]&rd_wr,DATAOUT);
	tristate32bit TSB22(DFF_OUT[22],DECODER_OUT[22]&rd_wr,DATAOUT);
	tristate32bit TSB23(DFF_OUT[23],DECODER_OUT[23]&rd_wr,DATAOUT);
	tristate32bit TSB24(DFF_OUT[24],DECODER_OUT[24]&rd_wr,DATAOUT);
	tristate32bit TSB25(DFF_OUT[25],DECODER_OUT[25]&rd_wr,DATAOUT);
	tristate32bit TSB26(DFF_OUT[26],DECODER_OUT[26]&rd_wr,DATAOUT);
	tristate32bit TSB27(DFF_OUT[27],DECODER_OUT[27]&rd_wr,DATAOUT);
	tristate32bit TSB28(DFF_OUT[28],DECODER_OUT[28]&rd_wr,DATAOUT);
	tristate32bit TSB29(DFF_OUT[29],DECODER_OUT[29]&rd_wr,DATAOUT);
	tristate32bit TSB30(DFF_OUT[30],DECODER_OUT[30]&rd_wr,DATAOUT);
	tristate32bit TSB31(DFF_OUT[31],DECODER_OUT[31]&rd_wr,DATAOUT);
	tristate32bit TSB32(DFF_OUT[32],DECODER_OUT[32]&rd_wr,DATAOUT);
	tristate32bit TSB33(DFF_OUT[33],DECODER_OUT[33]&rd_wr,DATAOUT);
	tristate32bit TSB34(DFF_OUT[34],DECODER_OUT[34]&rd_wr,DATAOUT);
	tristate32bit TSB35(DFF_OUT[35],DECODER_OUT[35]&rd_wr,DATAOUT);
	tristate32bit TSB36(DFF_OUT[36],DECODER_OUT[36]&rd_wr,DATAOUT);
	tristate32bit TSB37(DFF_OUT[37],DECODER_OUT[37]&rd_wr,DATAOUT);
	tristate32bit TSB38(DFF_OUT[38],DECODER_OUT[38]&rd_wr,DATAOUT);
	tristate32bit TSB39(DFF_OUT[39],DECODER_OUT[39]&rd_wr,DATAOUT);
	tristate32bit TSB40(DFF_OUT[40],DECODER_OUT[40]&rd_wr,DATAOUT);
	tristate32bit TSB41(DFF_OUT[41],DECODER_OUT[41]&rd_wr,DATAOUT);
	tristate32bit TSB42(DFF_OUT[42],DECODER_OUT[42]&rd_wr,DATAOUT);
	tristate32bit TSB43(DFF_OUT[43],DECODER_OUT[43]&rd_wr,DATAOUT);
	tristate32bit TSB44(DFF_OUT[44],DECODER_OUT[44]&rd_wr,DATAOUT);
	tristate32bit TSB45(DFF_OUT[45],DECODER_OUT[45]&rd_wr,DATAOUT);
	tristate32bit TSB46(DFF_OUT[46],DECODER_OUT[46]&rd_wr,DATAOUT);
	tristate32bit TSB47(DFF_OUT[47],DECODER_OUT[47]&rd_wr,DATAOUT);
	tristate32bit TSB48(DFF_OUT[48],DECODER_OUT[48]&rd_wr,DATAOUT);
	tristate32bit TSB49(DFF_OUT[49],DECODER_OUT[49]&rd_wr,DATAOUT);
	tristate32bit TSB50(DFF_OUT[50],DECODER_OUT[50]&rd_wr,DATAOUT);
	tristate32bit TSB51(DFF_OUT[51],DECODER_OUT[51]&rd_wr,DATAOUT);
	tristate32bit TSB52(DFF_OUT[52],DECODER_OUT[52]&rd_wr,DATAOUT);
	tristate32bit TSB53(DFF_OUT[53],DECODER_OUT[53]&rd_wr,DATAOUT);
	tristate32bit TSB54(DFF_OUT[54],DECODER_OUT[54]&rd_wr,DATAOUT);
	tristate32bit TSB55(DFF_OUT[55],DECODER_OUT[55]&rd_wr,DATAOUT);
	tristate32bit TSB56(DFF_OUT[56],DECODER_OUT[56]&rd_wr,DATAOUT);
	tristate32bit TSB57(DFF_OUT[57],DECODER_OUT[57]&rd_wr,DATAOUT);
	tristate32bit TSB58(DFF_OUT[58],DECODER_OUT[58]&rd_wr,DATAOUT);
	tristate32bit TSB59(DFF_OUT[59],DECODER_OUT[59]&rd_wr,DATAOUT);
	tristate32bit TSB60(DFF_OUT[60],DECODER_OUT[60]&rd_wr,DATAOUT);
	tristate32bit TSB61(DFF_OUT[61],DECODER_OUT[61]&rd_wr,DATAOUT);
	tristate32bit TSB62(DFF_OUT[62],DECODER_OUT[62]&rd_wr,DATAOUT);
	tristate32bit TSB63(DFF_OUT[63],DECODER_OUT[63]&rd_wr,DATAOUT);
	tristate32bit TSB64(DFF_OUT[64],DECODER_OUT[64]&rd_wr,DATAOUT);
	tristate32bit TSB65(DFF_OUT[65],DECODER_OUT[65]&rd_wr,DATAOUT);
	tristate32bit TSB66(DFF_OUT[66],DECODER_OUT[66]&rd_wr,DATAOUT);
	tristate32bit TSB67(DFF_OUT[67],DECODER_OUT[67]&rd_wr,DATAOUT);
	tristate32bit TSB68(DFF_OUT[68],DECODER_OUT[68]&rd_wr,DATAOUT);
	tristate32bit TSB69(DFF_OUT[69],DECODER_OUT[69]&rd_wr,DATAOUT);
	tristate32bit TSB70(DFF_OUT[70],DECODER_OUT[70]&rd_wr,DATAOUT);
	tristate32bit TSB71(DFF_OUT[71],DECODER_OUT[71]&rd_wr,DATAOUT);
	tristate32bit TSB72(DFF_OUT[72],DECODER_OUT[72]&rd_wr,DATAOUT);
	tristate32bit TSB73(DFF_OUT[73],DECODER_OUT[73]&rd_wr,DATAOUT);
	tristate32bit TSB74(DFF_OUT[74],DECODER_OUT[74]&rd_wr,DATAOUT);
	tristate32bit TSB75(DFF_OUT[75],DECODER_OUT[75]&rd_wr,DATAOUT);
	tristate32bit TSB76(DFF_OUT[76],DECODER_OUT[76]&rd_wr,DATAOUT);
	tristate32bit TSB77(DFF_OUT[77],DECODER_OUT[77]&rd_wr,DATAOUT);
	tristate32bit TSB78(DFF_OUT[78],DECODER_OUT[78]&rd_wr,DATAOUT);
	tristate32bit TSB79(DFF_OUT[79],DECODER_OUT[79]&rd_wr,DATAOUT);
	tristate32bit TSB80(DFF_OUT[80],DECODER_OUT[80]&rd_wr,DATAOUT);
	tristate32bit TSB81(DFF_OUT[81],DECODER_OUT[81]&rd_wr,DATAOUT);
	tristate32bit TSB82(DFF_OUT[82],DECODER_OUT[82]&rd_wr,DATAOUT);
	tristate32bit TSB83(DFF_OUT[83],DECODER_OUT[83]&rd_wr,DATAOUT);
	tristate32bit TSB84(DFF_OUT[84],DECODER_OUT[84]&rd_wr,DATAOUT);
	tristate32bit TSB85(DFF_OUT[85],DECODER_OUT[85]&rd_wr,DATAOUT);
	tristate32bit TSB86(DFF_OUT[86],DECODER_OUT[86]&rd_wr,DATAOUT);
	tristate32bit TSB87(DFF_OUT[87],DECODER_OUT[87]&rd_wr,DATAOUT);
	tristate32bit TSB88(DFF_OUT[88],DECODER_OUT[88]&rd_wr,DATAOUT);
	tristate32bit TSB89(DFF_OUT[89],DECODER_OUT[89]&rd_wr,DATAOUT);
	tristate32bit TSB90(DFF_OUT[90],DECODER_OUT[90]&rd_wr,DATAOUT);
	tristate32bit TSB91(DFF_OUT[91],DECODER_OUT[91]&rd_wr,DATAOUT);
	tristate32bit TSB92(DFF_OUT[92],DECODER_OUT[92]&rd_wr,DATAOUT);
	tristate32bit TSB93(DFF_OUT[93],DECODER_OUT[93]&rd_wr,DATAOUT);
	tristate32bit TSB94(DFF_OUT[94],DECODER_OUT[94]&rd_wr,DATAOUT);
	tristate32bit TSB95(DFF_OUT[95],DECODER_OUT[95]&rd_wr,DATAOUT);
	tristate32bit TSB96(DFF_OUT[96],DECODER_OUT[96]&rd_wr,DATAOUT);
	tristate32bit TSB97(DFF_OUT[97],DECODER_OUT[97]&rd_wr,DATAOUT);
	tristate32bit TSB98(DFF_OUT[98],DECODER_OUT[98]&rd_wr,DATAOUT);
	tristate32bit TSB99(DFF_OUT[99],DECODER_OUT[99]&rd_wr,DATAOUT);
	tristate32bit TSB100(DFF_OUT[100],DECODER_OUT[100]&rd_wr,DATAOUT);
	tristate32bit TSB101(DFF_OUT[101],DECODER_OUT[101]&rd_wr,DATAOUT);
	tristate32bit TSB102(DFF_OUT[102],DECODER_OUT[102]&rd_wr,DATAOUT);
	tristate32bit TSB103(DFF_OUT[103],DECODER_OUT[103]&rd_wr,DATAOUT);
	tristate32bit TSB104(DFF_OUT[104],DECODER_OUT[104]&rd_wr,DATAOUT);
	tristate32bit TSB105(DFF_OUT[105],DECODER_OUT[105]&rd_wr,DATAOUT);
	tristate32bit TSB106(DFF_OUT[106],DECODER_OUT[106]&rd_wr,DATAOUT);
	tristate32bit TSB107(DFF_OUT[107],DECODER_OUT[107]&rd_wr,DATAOUT);
	tristate32bit TSB108(DFF_OUT[108],DECODER_OUT[108]&rd_wr,DATAOUT);
	tristate32bit TSB109(DFF_OUT[109],DECODER_OUT[109]&rd_wr,DATAOUT);
	tristate32bit TSB110(DFF_OUT[110],DECODER_OUT[110]&rd_wr,DATAOUT);
	tristate32bit TSB111(DFF_OUT[111],DECODER_OUT[111]&rd_wr,DATAOUT);
	tristate32bit TSB112(DFF_OUT[112],DECODER_OUT[112]&rd_wr,DATAOUT);
	tristate32bit TSB113(DFF_OUT[113],DECODER_OUT[113]&rd_wr,DATAOUT);
	tristate32bit TSB114(DFF_OUT[114],DECODER_OUT[114]&rd_wr,DATAOUT);
	tristate32bit TSB115(DFF_OUT[115],DECODER_OUT[115]&rd_wr,DATAOUT);
	tristate32bit TSB116(DFF_OUT[116],DECODER_OUT[116]&rd_wr,DATAOUT);
	tristate32bit TSB117(DFF_OUT[117],DECODER_OUT[117]&rd_wr,DATAOUT);
	tristate32bit TSB118(DFF_OUT[118],DECODER_OUT[118]&rd_wr,DATAOUT);
	tristate32bit TSB119(DFF_OUT[119],DECODER_OUT[119]&rd_wr,DATAOUT);
	tristate32bit TSB120(DFF_OUT[120],DECODER_OUT[120]&rd_wr,DATAOUT);
	tristate32bit TSB121(DFF_OUT[121],DECODER_OUT[121]&rd_wr,DATAOUT);
	tristate32bit TSB122(DFF_OUT[122],DECODER_OUT[122]&rd_wr,DATAOUT);
	tristate32bit TSB123(DFF_OUT[123],DECODER_OUT[123]&rd_wr,DATAOUT);
	tristate32bit TSB124(DFF_OUT[124],DECODER_OUT[124]&rd_wr,DATAOUT);
	tristate32bit TSB125(DFF_OUT[125],DECODER_OUT[125]&rd_wr,DATAOUT);
	tristate32bit TSB126(DFF_OUT[126],DECODER_OUT[126]&rd_wr,DATAOUT);
	tristate32bit TSB127(DFF_OUT[127],DECODER_OUT[127]&rd_wr,DATAOUT);
	tristate32bit TSB128(DFF_OUT[128],DECODER_OUT[128]&rd_wr,DATAOUT);
	tristate32bit TSB129(DFF_OUT[129],DECODER_OUT[129]&rd_wr,DATAOUT);
	tristate32bit TSB130(DFF_OUT[130],DECODER_OUT[130]&rd_wr,DATAOUT);
	tristate32bit TSB131(DFF_OUT[131],DECODER_OUT[131]&rd_wr,DATAOUT);
	tristate32bit TSB132(DFF_OUT[132],DECODER_OUT[132]&rd_wr,DATAOUT);
	tristate32bit TSB133(DFF_OUT[133],DECODER_OUT[133]&rd_wr,DATAOUT);
	tristate32bit TSB134(DFF_OUT[134],DECODER_OUT[134]&rd_wr,DATAOUT);
	tristate32bit TSB135(DFF_OUT[135],DECODER_OUT[135]&rd_wr,DATAOUT);
	tristate32bit TSB136(DFF_OUT[136],DECODER_OUT[136]&rd_wr,DATAOUT);
	tristate32bit TSB137(DFF_OUT[137],DECODER_OUT[137]&rd_wr,DATAOUT);
	tristate32bit TSB138(DFF_OUT[138],DECODER_OUT[138]&rd_wr,DATAOUT);
	tristate32bit TSB139(DFF_OUT[139],DECODER_OUT[139]&rd_wr,DATAOUT);
	tristate32bit TSB140(DFF_OUT[140],DECODER_OUT[140]&rd_wr,DATAOUT);
	tristate32bit TSB141(DFF_OUT[141],DECODER_OUT[141]&rd_wr,DATAOUT);
	tristate32bit TSB142(DFF_OUT[142],DECODER_OUT[142]&rd_wr,DATAOUT);
	tristate32bit TSB143(DFF_OUT[143],DECODER_OUT[143]&rd_wr,DATAOUT);
	tristate32bit TSB144(DFF_OUT[144],DECODER_OUT[144]&rd_wr,DATAOUT);
	tristate32bit TSB145(DFF_OUT[145],DECODER_OUT[145]&rd_wr,DATAOUT);
	tristate32bit TSB146(DFF_OUT[146],DECODER_OUT[146]&rd_wr,DATAOUT);
	tristate32bit TSB147(DFF_OUT[147],DECODER_OUT[147]&rd_wr,DATAOUT);
	tristate32bit TSB148(DFF_OUT[148],DECODER_OUT[148]&rd_wr,DATAOUT);
	tristate32bit TSB149(DFF_OUT[149],DECODER_OUT[149]&rd_wr,DATAOUT);
	tristate32bit TSB150(DFF_OUT[150],DECODER_OUT[150]&rd_wr,DATAOUT);
	tristate32bit TSB151(DFF_OUT[151],DECODER_OUT[151]&rd_wr,DATAOUT);
	tristate32bit TSB152(DFF_OUT[152],DECODER_OUT[152]&rd_wr,DATAOUT);
	tristate32bit TSB153(DFF_OUT[153],DECODER_OUT[153]&rd_wr,DATAOUT);
	tristate32bit TSB154(DFF_OUT[154],DECODER_OUT[154]&rd_wr,DATAOUT);
	tristate32bit TSB155(DFF_OUT[155],DECODER_OUT[155]&rd_wr,DATAOUT);
	tristate32bit TSB156(DFF_OUT[156],DECODER_OUT[156]&rd_wr,DATAOUT);
	tristate32bit TSB157(DFF_OUT[157],DECODER_OUT[157]&rd_wr,DATAOUT);
	tristate32bit TSB158(DFF_OUT[158],DECODER_OUT[158]&rd_wr,DATAOUT);
	tristate32bit TSB159(DFF_OUT[159],DECODER_OUT[159]&rd_wr,DATAOUT);
	tristate32bit TSB160(DFF_OUT[160],DECODER_OUT[160]&rd_wr,DATAOUT);
	tristate32bit TSB161(DFF_OUT[161],DECODER_OUT[161]&rd_wr,DATAOUT);
	tristate32bit TSB162(DFF_OUT[162],DECODER_OUT[162]&rd_wr,DATAOUT);
	tristate32bit TSB163(DFF_OUT[163],DECODER_OUT[163]&rd_wr,DATAOUT);
	tristate32bit TSB164(DFF_OUT[164],DECODER_OUT[164]&rd_wr,DATAOUT);
	tristate32bit TSB165(DFF_OUT[165],DECODER_OUT[165]&rd_wr,DATAOUT);
	tristate32bit TSB166(DFF_OUT[166],DECODER_OUT[166]&rd_wr,DATAOUT);
	tristate32bit TSB167(DFF_OUT[167],DECODER_OUT[167]&rd_wr,DATAOUT);
	tristate32bit TSB168(DFF_OUT[168],DECODER_OUT[168]&rd_wr,DATAOUT);
	tristate32bit TSB169(DFF_OUT[169],DECODER_OUT[169]&rd_wr,DATAOUT);
	tristate32bit TSB170(DFF_OUT[170],DECODER_OUT[170]&rd_wr,DATAOUT);
	tristate32bit TSB171(DFF_OUT[171],DECODER_OUT[171]&rd_wr,DATAOUT);
	tristate32bit TSB172(DFF_OUT[172],DECODER_OUT[172]&rd_wr,DATAOUT);
	tristate32bit TSB173(DFF_OUT[173],DECODER_OUT[173]&rd_wr,DATAOUT);
	tristate32bit TSB174(DFF_OUT[174],DECODER_OUT[174]&rd_wr,DATAOUT);
	tristate32bit TSB175(DFF_OUT[175],DECODER_OUT[175]&rd_wr,DATAOUT);
	tristate32bit TSB176(DFF_OUT[176],DECODER_OUT[176]&rd_wr,DATAOUT);
	tristate32bit TSB177(DFF_OUT[177],DECODER_OUT[177]&rd_wr,DATAOUT);
	tristate32bit TSB178(DFF_OUT[178],DECODER_OUT[178]&rd_wr,DATAOUT);
	tristate32bit TSB179(DFF_OUT[179],DECODER_OUT[179]&rd_wr,DATAOUT);
	tristate32bit TSB180(DFF_OUT[180],DECODER_OUT[180]&rd_wr,DATAOUT);
	tristate32bit TSB181(DFF_OUT[181],DECODER_OUT[181]&rd_wr,DATAOUT);
	tristate32bit TSB182(DFF_OUT[182],DECODER_OUT[182]&rd_wr,DATAOUT);
	tristate32bit TSB183(DFF_OUT[183],DECODER_OUT[183]&rd_wr,DATAOUT);
	tristate32bit TSB184(DFF_OUT[184],DECODER_OUT[184]&rd_wr,DATAOUT);
	tristate32bit TSB185(DFF_OUT[185],DECODER_OUT[185]&rd_wr,DATAOUT);
	tristate32bit TSB186(DFF_OUT[186],DECODER_OUT[186]&rd_wr,DATAOUT);
	tristate32bit TSB187(DFF_OUT[187],DECODER_OUT[187]&rd_wr,DATAOUT);
	tristate32bit TSB188(DFF_OUT[188],DECODER_OUT[188]&rd_wr,DATAOUT);
	tristate32bit TSB189(DFF_OUT[189],DECODER_OUT[189]&rd_wr,DATAOUT);
	tristate32bit TSB190(DFF_OUT[190],DECODER_OUT[190]&rd_wr,DATAOUT);
	tristate32bit TSB191(DFF_OUT[191],DECODER_OUT[191]&rd_wr,DATAOUT);
	tristate32bit TSB192(DFF_OUT[192],DECODER_OUT[192]&rd_wr,DATAOUT);
	tristate32bit TSB193(DFF_OUT[193],DECODER_OUT[193]&rd_wr,DATAOUT);
	tristate32bit TSB194(DFF_OUT[194],DECODER_OUT[194]&rd_wr,DATAOUT);
	tristate32bit TSB195(DFF_OUT[195],DECODER_OUT[195]&rd_wr,DATAOUT);
	tristate32bit TSB196(DFF_OUT[196],DECODER_OUT[196]&rd_wr,DATAOUT);
	tristate32bit TSB197(DFF_OUT[197],DECODER_OUT[197]&rd_wr,DATAOUT);
	tristate32bit TSB198(DFF_OUT[198],DECODER_OUT[198]&rd_wr,DATAOUT);
	tristate32bit TSB199(DFF_OUT[199],DECODER_OUT[199]&rd_wr,DATAOUT);
	tristate32bit TSB200(DFF_OUT[200],DECODER_OUT[200]&rd_wr,DATAOUT);
	tristate32bit TSB201(DFF_OUT[201],DECODER_OUT[201]&rd_wr,DATAOUT);
	tristate32bit TSB202(DFF_OUT[202],DECODER_OUT[202]&rd_wr,DATAOUT);
	tristate32bit TSB203(DFF_OUT[203],DECODER_OUT[203]&rd_wr,DATAOUT);
	tristate32bit TSB204(DFF_OUT[204],DECODER_OUT[204]&rd_wr,DATAOUT);
	tristate32bit TSB205(DFF_OUT[205],DECODER_OUT[205]&rd_wr,DATAOUT);
	tristate32bit TSB206(DFF_OUT[206],DECODER_OUT[206]&rd_wr,DATAOUT);
	tristate32bit TSB207(DFF_OUT[207],DECODER_OUT[207]&rd_wr,DATAOUT);
	tristate32bit TSB208(DFF_OUT[208],DECODER_OUT[208]&rd_wr,DATAOUT);
	tristate32bit TSB209(DFF_OUT[209],DECODER_OUT[209]&rd_wr,DATAOUT);
	tristate32bit TSB210(DFF_OUT[210],DECODER_OUT[210]&rd_wr,DATAOUT);
	tristate32bit TSB211(DFF_OUT[211],DECODER_OUT[211]&rd_wr,DATAOUT);
	tristate32bit TSB212(DFF_OUT[212],DECODER_OUT[212]&rd_wr,DATAOUT);
	tristate32bit TSB213(DFF_OUT[213],DECODER_OUT[213]&rd_wr,DATAOUT);
	tristate32bit TSB214(DFF_OUT[214],DECODER_OUT[214]&rd_wr,DATAOUT);
	tristate32bit TSB215(DFF_OUT[215],DECODER_OUT[215]&rd_wr,DATAOUT);
	tristate32bit TSB216(DFF_OUT[216],DECODER_OUT[216]&rd_wr,DATAOUT);
	tristate32bit TSB217(DFF_OUT[217],DECODER_OUT[217]&rd_wr,DATAOUT);
	tristate32bit TSB218(DFF_OUT[218],DECODER_OUT[218]&rd_wr,DATAOUT);
	tristate32bit TSB219(DFF_OUT[219],DECODER_OUT[219]&rd_wr,DATAOUT);
	tristate32bit TSB220(DFF_OUT[220],DECODER_OUT[220]&rd_wr,DATAOUT);
	tristate32bit TSB221(DFF_OUT[221],DECODER_OUT[221]&rd_wr,DATAOUT);
	tristate32bit TSB222(DFF_OUT[222],DECODER_OUT[222]&rd_wr,DATAOUT);
	tristate32bit TSB223(DFF_OUT[223],DECODER_OUT[223]&rd_wr,DATAOUT);
	tristate32bit TSB224(DFF_OUT[224],DECODER_OUT[224]&rd_wr,DATAOUT);
	tristate32bit TSB225(DFF_OUT[225],DECODER_OUT[225]&rd_wr,DATAOUT);
	tristate32bit TSB226(DFF_OUT[226],DECODER_OUT[226]&rd_wr,DATAOUT);
	tristate32bit TSB227(DFF_OUT[227],DECODER_OUT[227]&rd_wr,DATAOUT);
	tristate32bit TSB228(DFF_OUT[228],DECODER_OUT[228]&rd_wr,DATAOUT);
	tristate32bit TSB229(DFF_OUT[229],DECODER_OUT[229]&rd_wr,DATAOUT);
	tristate32bit TSB230(DFF_OUT[230],DECODER_OUT[230]&rd_wr,DATAOUT);
	tristate32bit TSB231(DFF_OUT[231],DECODER_OUT[231]&rd_wr,DATAOUT);
	tristate32bit TSB232(DFF_OUT[232],DECODER_OUT[232]&rd_wr,DATAOUT);
	tristate32bit TSB233(DFF_OUT[233],DECODER_OUT[233]&rd_wr,DATAOUT);
	tristate32bit TSB234(DFF_OUT[234],DECODER_OUT[234]&rd_wr,DATAOUT);
	tristate32bit TSB235(DFF_OUT[235],DECODER_OUT[235]&rd_wr,DATAOUT);
	tristate32bit TSB236(DFF_OUT[236],DECODER_OUT[236]&rd_wr,DATAOUT);
	tristate32bit TSB237(DFF_OUT[237],DECODER_OUT[237]&rd_wr,DATAOUT);
	tristate32bit TSB238(DFF_OUT[238],DECODER_OUT[238]&rd_wr,DATAOUT);
	tristate32bit TSB239(DFF_OUT[239],DECODER_OUT[239]&rd_wr,DATAOUT);
	tristate32bit TSB240(DFF_OUT[240],DECODER_OUT[240]&rd_wr,DATAOUT);
	tristate32bit TSB241(DFF_OUT[241],DECODER_OUT[241]&rd_wr,DATAOUT);
	tristate32bit TSB242(DFF_OUT[242],DECODER_OUT[242]&rd_wr,DATAOUT);
	tristate32bit TSB243(DFF_OUT[243],DECODER_OUT[243]&rd_wr,DATAOUT);
	tristate32bit TSB244(DFF_OUT[244],DECODER_OUT[244]&rd_wr,DATAOUT);
	tristate32bit TSB245(DFF_OUT[245],DECODER_OUT[245]&rd_wr,DATAOUT);
	tristate32bit TSB246(DFF_OUT[246],DECODER_OUT[246]&rd_wr,DATAOUT);
	tristate32bit TSB247(DFF_OUT[247],DECODER_OUT[247]&rd_wr,DATAOUT);
	tristate32bit TSB248(DFF_OUT[248],DECODER_OUT[248]&rd_wr,DATAOUT);
	tristate32bit TSB249(DFF_OUT[249],DECODER_OUT[249]&rd_wr,DATAOUT);
	tristate32bit TSB250(DFF_OUT[250],DECODER_OUT[250]&rd_wr,DATAOUT);
	tristate32bit TSB251(DFF_OUT[251],DECODER_OUT[251]&rd_wr,DATAOUT);
	tristate32bit TSB252(DFF_OUT[252],DECODER_OUT[252]&rd_wr,DATAOUT);
	tristate32bit TSB253(DFF_OUT[253],DECODER_OUT[253]&rd_wr,DATAOUT);
	tristate32bit TSB254(DFF_OUT[254],DECODER_OUT[254]&rd_wr,DATAOUT);
	tristate32bit TSB255(DFF_OUT[255],DECODER_OUT[255]&rd_wr,DATAOUT);
	
endmodule

`endif
